-----------------------------------------------------------------
-- (c) Copyright 2017
-- Critical Software S.A.
-- All Rights Reserved
-----------------------------------------------------------------
-- Project     : VCU
-- Filename    : TC_RS088_183
-- Module      : VCU Timing System
-- Revision    : 1.0
-- Date        : 30 Jan 2020
-- Author      : CABelchior
-----------------------------------------------------------------
-- Description : Check that all minor error status flags shall be reported to the following external means
-----------------------------------------------------------------
-- Requirements:
--    FPGA-REQ-88
--    FPGA-REQ-183
-----------------------------------------------------------------
-- History:
-- Revision 1.0 - 30 Jan 2020
--    - CABelchior (2.0): CCN04 Updates (also test bench updates)
-----------------------------------------------------------------
-- Notes:
--
-- sim -tc TC_RS088_183 -numstdoff -nocov
-- log -r /*
--
-- 88    All minor error status flags shall be reported to the following external means:
--       - TMS
--       - LED Display
--
-- 183   (...) The display minor fault and major fault pins should be driven high when their 
--       respective faults are found.
--
--   Minor Fault IF - Inputs
--   -----------------------
--   input_flt_i => (input_if::fault_o)
--   spd_urng_i  => (input_if::spd_urng_o)
--   spd_orng_i  => (input_if::spd_orng_o)
--   spd_err_i   => (input_if::spd_err_o)
--   dry_flt_i   => (output_if::dry_flt_o)
--   wet_flt_i   => (output_if::wet_flt_o)
--
--   fault_o <= st_fault_s                        - FPGA-REQ-188
--              OR (pwm0_fault_s OR pwm1_fault_s) - FPGA-REQ-36
--              OR OR_REDUCE(compare_fault_s)     - FPGA-REQ-22
--              OR (ps1_fail_s1 OR ps2_fail_s1)   - FPGA-REQ-201
--
--   spd_urng_o                                   - FPGA-REQ-202
--
--   spd_orng_o                                   - FPGA-REQ-202
--
--   spd_err_o                                    - FPGA-REQ-202
--
--   dry_flt_o                                    - FPGA-REQ-67
--
--   wet_flt_o                                    - FPGA-REQ-66
--
-- Aditional notes: 
-- ----------------------
-- As stated in ARCHITECTURE DESIGN AND INTERFACE SPECIFICATION document, the Minor Fault block 
-- aggregates all inputs that contribute to the generation of this fault type. The output of this 
-- block is simply an OR of all its inputs.
-- 
-- The input_flt_i signal is an input from the Input IF HLB, specifically from the Fault Calc block 
-- described in section 3.4.2.2. 
--
-- The spd_urng_i, spd_orng_i and spd_err_i signals correspond to the analog speed under-range, 
-- over-range and reading faults processed by the Analog IF block within the Input IF HLB described 
-- in Section 3.4.2.8.
--
-- Finally, the dry_flt_i and wet_flt_i vectors are the faults generated by the Output IF block, 
-- described in section, 3.4.7 for all outputs that fail the feedback comparison routine according 
-- to [RD-2] section 4.2.
--
-- Aditional notes: 
-- ----------------------
-- minor_flt_report_s         <= tms_minor_fault_o AND disp_minor_fault_o;
-- major_flt_report_s         <= tms_major_fault_o AND disp_major_fault_o;
-----------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.All;
USE IEEE.NUMERIC_STD.All;
USE IEEE.MATH_REAL.All;

LIBRARY modelsim_lib;
USE     modelsim_lib.util.ALL;
USE WORK.testify_p.ALL;

ARCHITECTURE TC_RS088_183 OF hcmt_cpld_tc_top IS

   --------------------------------------------------------
   -- Applicable Constants
   --------------------------------------------------------

   --------------------------------------------------------
   -- Spy Probes
   --------------------------------------------------------

   --------------------------------------------------------
   -- User Signals
   --------------------------------------------------------
   SIGNAL s_usr_sigout_s                          : tfy_user_out;
   SIGNAL s_usr_sigin_s                           : tfy_user_in;
   SIGNAL pwm_func_model_data_s                   : pwm_func_model_inputs := C_PWM_FUNC_MODEL_INPUTS_INIT;   
   SIGNAL st_ch1_in_ctrl_s                        : ST_BEHAVIOR_CH1;
   SIGNAL st_ch2_in_ctrl_s                        : ST_BEHAVIOR_CH2;

   SIGNAL minor_flt_report_s                      : STD_LOGIC := '0';

BEGIN

   p_steps: PROCESS

      --------------------------------------------------------
      -- Common Test Case variable declarations
      --------------------------------------------------------
      VARIABLE pass                              : BOOLEAN := true;

      --------------------------------------------------------
      -- Other Testcase Variables
      --------------------------------------------------------
      VARIABLE ta, tb, tc, td, te, tf, tg        : TIME;
      VARIABLE dt                                : TIME;

      --------------------------------------------------------
      -- Procedures & Functions
      --------------------------------------------------------

      PROCEDURE Set_Speed_Cases(spd_cases : NATURAL) IS
      BEGIN
         uut_in.spd_over_spd_s     <= C_SPEED_VALUES(spd_cases)(7);
         uut_in.spd_h110kmh_s      <= C_SPEED_VALUES(spd_cases)(6);
         uut_in.spd_h90kmh_s       <= C_SPEED_VALUES(spd_cases)(5);
         uut_in.spd_h75kmh_s       <= C_SPEED_VALUES(spd_cases)(4);
         uut_in.spd_h25kmh_a_s     <= C_SPEED_VALUES(spd_cases)(3);
         uut_in.spd_h25kmh_b_s     <= C_SPEED_VALUES(spd_cases)(3);
         uut_in.spd_h23kmh_a_s     <= C_SPEED_VALUES(spd_cases)(2);
         uut_in.spd_h23kmh_b_s     <= C_SPEED_VALUES(spd_cases)(2);
         uut_in.spd_h3kmh_s        <= C_SPEED_VALUES(spd_cases)(1);
         uut_in.spd_l3kmh_s        <= C_SPEED_VALUES(spd_cases)(0);
      END PROCEDURE Set_Speed_Cases;

      PROCEDURE Reset_UUT (Step : STRING) IS 
      BEGIN
         -------------------------------------------------
         tfy_wr_step( report_file, now, Step, 
            "Configure and reset UUT to clear all persistent errors");

         -------------------------------------------------
         tfy_wr_step( report_file, now, Step & ".1", 
            "Configure all functional models to normal behavior");
         st_ch1_in_ctrl_s        <= (OTHERS => C_ST_FUNC_MODEL_ARRAY_INIT);
         st_ch2_in_ctrl_s        <= (OTHERS => C_ST_FUNC_MODEL_ARRAY_INIT);
         fb_func_model_behaviour <= C_OUT_FB_FUNC_MODEL_BEHAVIOUR_INIT;
         pwm_func_model_data_s   <= C_PWM_FUNC_MODEL_INPUTS_INIT;

         -------------------------------------------------
         tfy_wr_step( report_file, now, Step & ".2", 
            "Set all dual channel inputs to '0'");
         uut_in.vigi_pb_ch1_s          <= '0';
         uut_in.vigi_pb_ch2_s          <= '0';
   
         uut_in.zero_spd_ch1_s         <= '0';
         uut_in.zero_spd_ch2_s         <= '0';
         
         uut_in.hcs_mode_ch1_s         <= '0';
         uut_in.hcs_mode_ch2_s         <= '0';
         
         uut_in.bcp_75_ch1_s           <= '0';
         uut_in.bcp_75_ch2_s           <= '0';
         
         uut_in.not_isol_ch1_s         <= '0';
         uut_in.not_isol_ch2_s         <= '0';
         
         uut_in.cab_act_ch1_s          <= '0';
         uut_in.cab_act_ch2_s          <= '0';
         
         uut_in.spd_lim_override_ch1_s <= '0';
         uut_in.spd_lim_override_ch2_s <= '0';
         
         uut_in.driverless_ch1_s       <= '0';
         uut_in.driverless_ch2_s       <= '0';
         
         uut_in.spd_lim_ch1_s          <= '0';
         uut_in.spd_lim_ch2_s          <= '0';

         -------------------------------------------------
         tfy_wr_step( report_file, now, Step & ".3", 
            "Set all single channel inputs to '0'");
         uut_in.horn_low_s             <= '0';
         uut_in.horn_high_s            <= '0';
         uut_in.hl_low_s               <= '0';
         uut_in.w_wiper_pb_s           <= '0';
         uut_in.ss_bypass_pb_s         <= '0';

         -------------------------------------------------
         tfy_wr_step( report_file, now, Step & ".4", 
            "Set all feedback inputs for digital outputs to 'Z'");
         uut_in.light_out_fb_s               <= 'Z';

         uut_in.tms_pb_fb_s                  <= 'Z';
         uut_in.tms_spd_lim_overridden_fb_s  <= 'Z';
         uut_in.tms_rst_fb_s                 <= 'Z';
         uut_in.tms_penalty_stat_fb_s        <= 'Z';
         uut_in.tms_major_fault_fb_s         <= 'Z';
         uut_in.tms_minor_fault_fb_s         <= 'Z';
         uut_in.tms_depressed_fb_s           <= 'Z';
         uut_in.tms_suppressed_fb_s          <= 'Z';
         uut_in.tms_vis_warn_stat_fb_s       <= 'Z';
         uut_in.tms_spd_lim_stat_fb_s        <= 'Z';
      
         uut_in.buzzer_out_fb_s              <= 'Z';
      
         uut_in.penalty2_fb_s                <= 'Z';
         uut_in.penalty1_fb_s                <= 'Z';
         uut_in.rly_fb3_3V_s                 <= 'Z';
         uut_in.rly_fb2_3V_s                 <= 'Z';
         uut_in.rly_fb1_3V_s                 <= 'Z';

         -------------------------------------------------
         tfy_wr_step( report_file, now, Step & ".5", 
            "Set analog speed to [0 - 3 km/h]");
         Set_Speed_Cases(1);               -- Analog Speed -> 0 – 3 km/h

         -------------------------------------------------
         tfy_wr_step( report_file, now, Step & ".6", 
            "Set power supply 1&2 failure status to '1', i.e. OK");
         uut_in.ps1_stat_s        <= '1';  -- Power supply 1 Status OK
         uut_in.ps2_stat_s        <= '1';  -- Power supply 1 Status OK

         -------------------------------------------------
         tfy_wr_step( report_file, now, Step & ".7", 
            "Set CH1 and CH2 external self-test circuitry signal to '0'");
         uut_in.force_fault_ch1_s <= '0';  -- External CH1 self-test circuitry OK
         uut_in.force_fault_ch2_s <= '0';  -- External CH2 self-test circuitry OK

         -------------------------------------------------
         tfy_wr_step( report_file, now, Step & ".8", 
            "Reset UUT and wait for 10ms for system power-up");
         uut_in.arst_n_s     <= '0';       -- Reset UUT
         wait_for_clk_cycles(30, Clk);
         uut_in.arst_n_s     <= '1';
         WAIT FOR 10 ms;                   -- System Power Up

      END PROCEDURE Reset_UUT;

   BEGIN

      --------------------------------------------------------
      -- Testcase Start Sequence
      --------------------------------------------------------
      tfy_tc_start(
         report_fname   => "TC_RS088_183.rep",
         report_file    => report_file,
         project_name   => "VCU",
         tc_name        => "TC_RS088_183",
         test_module    => "VCU Timing System",
         tc_revision    => "1.0",
         tc_date        => "30 Jan 2020",
         tester_name    => "CABelchior",
         tc_description => "Check that all minor error status flags shall be reported to the following external means",
         tb_name        => "hcmt_cpld_top_tb",
         dut_name       => "hcmt_cpld_top_tb",
         s_usr_sigin_s  => s_usr_sigin_s,
         s_usr_sigout_s => s_usr_sigout_s
      );   

      --------------------------------------------------------
      -- Link Spy Probes
      --------------------------------------------------------

      --------------------------------------------------------
      -- Link Drive Probes
      --------------------------------------------------------

      --------------------------------------------------------
      -- Initializations
      --------------------------------------------------------
      tfy_wr_console(" [*] Simulation Init");
      uut_in                   <= f_uutinit('Z');
      uut_inout.SDAInout       <= 'Z';
      uut_in.arst_n_s          <= '0';
      s_usr_sigin_s.bfm_pass   <= TRUE;

      --------------------------------------------------------
      -- Testcase Steps
      --------------------------------------------------------

      --==============
      -- Step 1
      --==============

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_console(" [*] Step 1: -------------------------------------------#");
      tfy_wr_step( report_file, now, "1",
         "The specification of Minor Fault generation due to signal 'input_flt_i' is done at:");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "1.1",
         "FPGA-REQ-188 - Any fault reported by the Self-Test routine");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "1.1.1",
         "The verification of this statement occurs at: TC_RS016_023_027_012_188");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "1.2",
         "FPGA-REQ-36 - Any condition causing either or both PWM being masked permanently");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "1.2.1",
         "The verification of this statement occurs at: TC_RS036_191_192_084_194");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "1.3",
         "FPGA-REQ-22 - If there is a fault at any dual channel signal comparison for a sufficient time to be considered permanent");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "1.3.1",
         "The verification of this statement occurs at: TC_RS018_019_020_021_022_203");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "1.4",
         "FPGA-REQ-201 - If either the power supply 1 or 2 status signals are low for a sufficient time to be considered a permanent fault");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "1.4.1",
         "The verification of this statement occurs at: TC_RS201");


      --==============
      -- Step 2
      --==============

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_console(" [*] Step 2: -------------------------------------------#");
      tfy_wr_step( report_file, now, "2",
         "The specification of Minor Fault generation due to signal 'spd_urng_i' is done at:");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "2.1",
         "FPGA-REQ-202 - If the speed value indicates an error of type 'Under Range' for a sufficient time to be considered a permanent fault");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "2.1.1",
         "The verification of this statement occurs at: TC_RS040_041_042_043_202_179");


      --==============
      -- Step 3
      --==============

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_console(" [*] Step 3: -------------------------------------------#");
      tfy_wr_step( report_file, now, "3",
         "The specification of Minor Fault generation due to signal 'spd_orng_i' is done at:");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "3.1",
         "FPGA-REQ-202 - If the speed value indicates an error of type 'Over Range' for a sufficient time to be considered a permanent fault");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "3.1.1",
         "The verification of this statement occurs at: TC_RS040_041_042_043_202_179");


      --==============
      -- Step 4
      --==============

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_console(" [*] Step 4: -------------------------------------------#");
      tfy_wr_step( report_file, now, "4",
         "The specification of Minor Fault generation due to signal 'spd_err_i' is done at:");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "4.1",
         "FPGA-REQ-202 - If the speed value indicates an error of type 'Invalid Speed' for a sufficient time to be considered a permanent fault");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "4.1.1",
         "The verification of this statement occurs at: TC_RS040_041_042_043_202_179");


      --==============
      -- Step 5
      --==============

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_console(" [*] Step 5: -------------------------------------------#");
      tfy_wr_step( report_file, now, "5",
         "The specification of Minor Fault generation due to signal 'dry_flt_i' is done at:");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "5.1",
         "FPGA-REQ-67 - If there is a fault at a dry output comparison for a sufficient time to be considered permanent");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "5.1.1",
         "The verification of this statement occurs at: TC_RS065_067_137_164");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "5.1.2",
         "The verification of this statement occurs at: TC_RS065_067_137_168");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "5.1.3",
         "The verification of this statement occurs at: TC_RS065_067_137_170");

         
      --==============
      -- Step 6
      --==============

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_console(" [*] Step 6: -------------------------------------------#");
      tfy_wr_step( report_file, now, "6",
         "The specification of Minor Fault generation due to signal 'wet_flt_i' is done at:");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "6.1",
         "FPGA-REQ-66 - If there is a fault at a wet output comparison for a sufficient time to be considered permanent");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "6.1.1",
         "The verification of this statement occurs at: TC_RS065_066_137_141");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "6.1.2",
         "The verification of this statement occurs at: TC_RS065_066_137_143");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "6.1.3",
         "The verification of this statement occurs at: TC_RS065_066_137_145");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "6.1.4",
         "The verification of this statement occurs at: TC_RS065_066_137_149");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "6.1.5",
         "The verification of this statement occurs at: TC_RS065_066_137_152");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "6.1.6",
         "The verification of this statement occurs at: TC_RS065_066_137_154");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "6.1.7",
         "The verification of this statement occurs at: TC_RS065_066_137_156");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "6.1.8",
         "The verification of this statement occurs at: TC_RS065_066_137_158");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "6.1.9",
         "The verification of this statement occurs at: TC_RS065_066_137_160");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "6.1.10",
         "The verification of this statement occurs at: TC_RS065_066_137_197");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "6.1.11",
         "The verification of this statement occurs at: TC_RS065_066_137_199");

      -----------------------------------------------------------------------------------------------------------
      tfy_wr_step( report_file, now, "6.1.12",
         "The verification of this statement occurs at: TC_RS065_066_137_212");

      --------------------------------------------------------
      -- END
      --------------------------------------------------------
      WAIT FOR 20 ms;
      --------------------------------------------------------
      -- Testcase End Sequence
      --------------------------------------------------------

      tfy_tc_end(
         tc_pass        => pass,
         report_file    => report_file,
         tc_name        => "TC_RS088_183",
         tb_name        => "hcmt_cpld_top_tb",
         dut_name       => "hcmt_cpld_tc_top",
         tester_name    => "CABelchior",
         tc_date        => "30 Jan 2020",
         s_usr_sigin_s  => s_usr_sigin_s,
         s_usr_sigout_s => s_usr_sigout_s    
      );

   END PROCESS p_steps;

   s_usr_sigin_s.test_select  <= test_select;
   s_usr_sigin_s.clk          <= Clk;
   test_done                  <= s_usr_sigout_s.test_done;
   pwm_func_model_data        <= pwm_func_model_data_s;
   st_ch1_in_ctrl_o           <= st_ch1_in_ctrl_s; 
   st_ch2_in_ctrl_o           <= st_ch2_in_ctrl_s; 
   
   minor_flt_report_s         <= uut_out.tms_minor_fault_s AND uut_out.disp_minor_fault_s;
END ARCHITECTURE TC_RS088_183;
